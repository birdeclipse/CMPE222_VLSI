magic
tech scmos
timestamp 1460581730
use INVX8  INVX8_3
timestamp 1460491589
transform 1 0 -16 0 -1 77
box -28 -58 10 25
use INVX8  INVX8_1
timestamp 1460491589
transform 1 0 4 0 -1 77
box -28 -58 10 25
use INVX8  INVX8_2
timestamp 1460491589
transform 1 0 24 0 -1 77
box -28 -58 10 25
use INVX8  INVX8_5
timestamp 1460491589
transform 1 0 -16 0 1 39
box -28 -58 10 25
use INVX8  INVX8_0
timestamp 1460491589
transform 1 0 4 0 1 39
box -28 -58 10 25
use INVX8  INVX8_4
timestamp 1460491589
transform 1 0 24 0 1 39
box -28 -58 10 25
use INVX8  INVX8_6
timestamp 1460491589
transform 1 0 -16 0 -1 -67
box -28 -58 10 25
use INVX8  INVX8_7
timestamp 1460491589
transform 1 0 4 0 -1 -67
box -28 -58 10 25
use INVX8  INVX8_8
timestamp 1460491589
transform 1 0 24 0 -1 -67
box -28 -58 10 25
<< end >>
