magic
tech scmos
timestamp 1460174537
<< nwell >>
rect -28 -9 10 25
<< pwell >>
rect -28 -40 11 -12
<< ntransistor >>
rect -10 -26 -8 -18
<< ptransistor >>
rect -10 -3 -8 13
<< ndiffusion >>
rect -11 -26 -10 -18
rect -8 -26 -7 -18
<< pdiffusion >>
rect -11 -3 -10 13
rect -8 -3 -7 13
<< ndcontact >>
rect -15 -26 -11 -18
rect -7 -26 -3 -18
<< pdcontact >>
rect -15 -3 -11 13
rect -7 -3 -3 13
<< psubstratepcontact >>
rect -20 -34 -16 -30
rect -2 -34 2 -30
<< nsubstratencontact >>
rect -20 17 -16 21
rect -2 17 2 21
<< polysilicon >>
rect -10 13 -8 15
rect -10 -7 -8 -3
rect -17 -11 -8 -7
rect -10 -18 -8 -11
rect -10 -28 -8 -26
<< polycontact >>
rect -21 -11 -17 -7
<< metal1 >>
rect -22 21 4 22
rect -22 17 -20 21
rect -16 17 -2 21
rect 2 17 4 21
rect -22 16 4 17
rect -15 13 -11 16
rect -7 -18 -3 -3
rect -15 -29 -11 -26
rect -22 -30 4 -29
rect -22 -34 -20 -30
rect -16 -34 -2 -30
rect 2 -34 4 -30
rect -22 -35 4 -34
<< metal2 >>
rect -25 -11 -17 -7
<< labels >>
rlabel metal2 -25 -11 -25 -11 3 +IN
rlabel nsubstratencontact -18 19 -18 19 1 +VDD
rlabel psubstratepcontact -18 -32 -18 -32 1 GND
<< end >>
