magic
tech scmos
timestamp 1460241879
use INVX8  INVX8_5
timestamp 1460237164
transform -1 0 -32 0 -1 69
box -28 -40 10 25
use INVX8  INVX8_0
timestamp 1460237164
transform -1 0 -8 0 -1 69
box -28 -40 10 25
use INVX8  INVX8_4
timestamp 1460237164
transform 1 0 35 0 -1 69
box -28 -40 10 25
use INVX8  INVX8_2
timestamp 1460237164
transform 1 0 -14 0 1 31
box -28 -40 10 25
use NAND2X2  NAND2X2_0
timestamp 1460241041
transform 1 0 7 0 1 9
box -25 -18 13 47
use INVX8  INVX8_1
timestamp 1460237164
transform 1 0 35 0 1 31
box -28 -40 10 25
use INVX8  INVX8_7
timestamp 1460237164
transform 1 0 -14 0 -1 -33
box -28 -40 10 25
use INVX8  INVX8_3
timestamp 1460237164
transform -1 0 -6 0 -1 -33
box -28 -40 10 25
use INVX8  INVX8_6
timestamp 1460237164
transform 1 0 35 0 -1 -33
box -28 -40 10 25
<< end >>
