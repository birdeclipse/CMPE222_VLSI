magic
tech scmos
timestamp 1460443535
<< nwell >>
rect -28 -9 10 25
<< pwell >>
rect -28 -40 10 -12
<< ntransistor >>
rect -10 -29 -8 -21
<< ptransistor >>
rect -10 -3 -8 13
<< ndiffusion >>
rect -11 -29 -10 -21
rect -8 -29 -7 -21
<< pdiffusion >>
rect -11 -3 -10 13
rect -8 -3 -7 13
<< ndcontact >>
rect -15 -29 -11 -21
rect -7 -29 -3 -21
<< pdcontact >>
rect -15 -3 -11 13
rect -7 -3 -3 13
<< psubstratepcontact >>
rect -21 -37 -17 -33
rect -1 -37 3 -33
<< nsubstratencontact >>
rect -21 17 -17 21
rect -1 17 3 21
<< polysilicon >>
rect -10 13 -8 15
rect -10 -8 -8 -3
rect -12 -12 -8 -8
rect -10 -21 -8 -12
rect -10 -31 -8 -29
<< polycontact >>
rect -16 -12 -12 -8
<< metal1 >>
rect -24 21 6 22
rect -24 17 -21 21
rect -17 17 -1 21
rect 3 17 6 21
rect -24 16 6 17
rect -15 13 -11 16
rect -16 -8 -12 -6
rect -7 -21 -3 -3
rect -15 -32 -11 -29
rect -24 -33 6 -32
rect -24 -37 -21 -33
rect -17 -37 -1 -33
rect 3 -37 6 -33
rect -24 -38 6 -37
<< labels >>
rlabel polycontact -14 -10 -14 -10 1 A
rlabel metal1 -5 -10 -5 -10 1 Z
rlabel nsubstratencontact -19 19 -19 19 1 +VDD
rlabel nsubstratencontact 1 19 1 19 1 +VDD
rlabel psubstratepcontact -19 -35 -19 -35 1 GND
rlabel psubstratepcontact 1 -35 1 -35 1 GND
<< end >>
