magic
tech scmos
timestamp 1460174745
use INVX8  INVX8_0
timestamp 1460174537
transform -1 0 -26 0 -1 53
box -28 -40 11 25
use NAND2X2  NAND2X2_0
timestamp 1460174587
transform 1 0 -11 0 1 4
box -25 -17 13 38
<< end >>
