magic
tech scmos
timestamp 1460150708
<< nwell >>
rect -35 0 -5 41
<< ntransistor >>
rect -21 -15 -19 -6
<< ptransistor >>
rect -21 8 -19 28
<< ndiffusion >>
rect -22 -15 -21 -6
rect -19 -15 -18 -6
<< pdiffusion >>
rect -22 8 -21 28
rect -19 8 -18 28
<< ndcontact >>
rect -26 -15 -22 -6
rect -18 -15 -14 -6
<< pdcontact >>
rect -26 8 -22 28
rect -18 8 -14 28
<< psubstratepcontact >>
rect -29 -26 -25 -22
rect -13 -26 -9 -22
<< nsubstratencontact >>
rect -29 33 -25 37
rect -14 33 -10 37
<< polysilicon >>
rect -21 28 -19 31
rect -21 3 -19 8
rect -25 -1 -19 3
rect -21 -6 -19 -1
rect -21 -20 -19 -15
<< polycontact >>
rect -29 -1 -25 3
<< metal1 >>
rect -32 37 -7 38
rect -32 33 -29 37
rect -25 33 -14 37
rect -10 33 -7 37
rect -32 32 -7 33
rect -26 28 -22 32
rect -33 -1 -29 3
rect -18 -6 -14 8
rect -26 -21 -22 -15
rect -32 -22 -6 -21
rect -32 -26 -29 -22
rect -25 -26 -13 -22
rect -9 -26 -6 -22
rect -32 -27 -6 -26
<< labels >>
rlabel metal1 -33 -1 -33 -1 3 in
rlabel metal1 -25 33 -25 33 1 vdd
rlabel metal1 -16 4 -16 4 1 out
rlabel metal1 -25 -26 -25 -26 1 gnd+
<< end >>
