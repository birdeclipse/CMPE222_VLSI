magic
tech scmos
timestamp 1460237164
<< nwell >>
rect -28 -9 10 25
<< pwell >>
rect -28 -40 10 -12
<< ntransistor >>
rect -10 -26 -8 -18
<< ptransistor >>
rect -10 -3 -8 13
<< ndiffusion >>
rect -11 -26 -10 -18
rect -8 -26 -7 -18
<< pdiffusion >>
rect -11 -3 -10 13
rect -8 -3 -7 13
<< ndcontact >>
rect -15 -26 -11 -18
rect -7 -26 -3 -18
<< pdcontact >>
rect -15 -3 -11 13
rect -7 -3 -3 13
<< psubstratepcontact >>
rect -11 -34 -7 -30
<< nsubstratencontact >>
rect -11 17 -7 21
<< polysilicon >>
rect -10 13 -8 15
rect -10 -18 -8 -3
rect -10 -28 -8 -26
<< polycontact >>
rect -14 -11 -10 -7
rect -3 -11 1 -7
<< metal1 >>
rect -22 21 4 22
rect -22 17 -11 21
rect -7 17 4 21
rect -22 16 4 17
rect -15 13 -11 16
rect -7 -18 -3 -3
rect -15 -29 -11 -26
rect -22 -30 4 -29
rect -22 -34 -11 -30
rect -7 -34 4 -30
rect -22 -35 4 -34
<< metal2 >>
rect -14 -11 -10 -7
rect -3 -11 1 -7
<< labels >>
rlabel nsubstratencontact -9 19 -9 19 1 +VDD
rlabel psubstratepcontact -9 -32 -9 -32 1 GND
rlabel polycontact -1 -9 -1 -9 1 OUT
rlabel metal2 -12 -9 -12 -9 1 IN
<< end >>
