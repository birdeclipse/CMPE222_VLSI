magic
tech scmos
timestamp 1460491589
<< nwell >>
rect -28 -9 10 25
<< pwell >>
rect -28 -58 10 -30
<< ntransistor >>
rect -10 -47 -8 -39
<< ptransistor >>
rect -10 -3 -8 13
<< ndiffusion >>
rect -11 -47 -10 -39
rect -8 -47 -7 -39
<< pdiffusion >>
rect -11 -3 -10 13
rect -8 -3 -7 13
<< ndcontact >>
rect -15 -47 -11 -39
rect -7 -47 -3 -39
<< pdcontact >>
rect -15 -3 -11 13
rect -7 -3 -3 13
<< psubstratepcontact >>
rect -21 -55 -17 -51
rect -1 -55 3 -51
<< nsubstratencontact >>
rect -21 17 -17 21
rect -1 17 3 21
<< polysilicon >>
rect -10 13 -8 15
rect -10 -39 -8 -3
rect -10 -49 -8 -47
<< polycontact >>
rect -14 -18 -10 -14
<< metal1 >>
rect -24 21 6 22
rect -24 17 -21 21
rect -17 17 -1 21
rect 3 17 6 21
rect -24 16 6 17
rect -15 13 -11 16
rect -7 -39 -3 -3
rect -15 -50 -11 -47
rect -24 -51 6 -50
rect -24 -55 -21 -51
rect -17 -55 -1 -51
rect 3 -55 6 -51
rect -24 -56 6 -55
<< labels >>
rlabel nsubstratencontact -19 19 -19 19 1 +VDD
rlabel nsubstratencontact 1 19 1 19 1 +VDD
rlabel psubstratepcontact -19 -53 -19 -53 1 GND
rlabel psubstratepcontact 1 -53 1 -53 1 GND
rlabel polycontact -12 -16 -12 -16 1 A
rlabel metal1 -5 -16 -5 -16 1 Z
<< end >>
