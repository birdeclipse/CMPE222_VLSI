magic
tech scmos
timestamp 1460444133
use NAND2X2  NAND2X2_5
timestamp 1460443965
transform 1 0 -48 0 -1 68
box -25 -18 13 47
use NAND2X2  NAND2X2_3
timestamp 1460443965
transform 1 0 -20 0 -1 68
box -25 -18 13 47
use NAND2X2  NAND2X2_4
timestamp 1460443965
transform 1 0 8 0 -1 68
box -25 -18 13 47
use NAND2X2  NAND2X2_2
timestamp 1460443965
transform 1 0 -48 0 1 -14
box -25 -18 13 47
use NAND2X2  NAND2X2_0
timestamp 1460443965
transform 1 0 -20 0 1 -14
box -25 -18 13 47
use NAND2X2  NAND2X2_1
timestamp 1460443965
transform 1 0 8 0 1 -14
box -25 -18 13 47
use NAND2X2  NAND2X2_6
timestamp 1460443965
transform 1 0 -48 0 -1 -40
box -25 -18 13 47
use NAND2X2  NAND2X2_7
timestamp 1460443965
transform 1 0 -20 0 -1 -40
box -25 -18 13 47
use NAND2X2  NAND2X2_8
timestamp 1460443965
transform 1 0 8 0 -1 -40
box -25 -18 13 47
<< end >>
