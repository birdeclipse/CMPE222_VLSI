magic
tech scmos
timestamp 1460443965
<< nwell >>
rect -25 13 13 47
<< pwell >>
rect -25 -18 13 10
<< ntransistor >>
rect -11 -7 -9 -3
rect -3 -7 -1 -3
<< ptransistor >>
rect -11 31 -9 35
rect -3 31 -1 35
<< ndiffusion >>
rect -12 -7 -11 -3
rect -9 -7 -3 -3
rect -1 -7 0 -3
<< pdiffusion >>
rect -12 31 -11 35
rect -9 31 -8 35
rect -4 31 -3 35
rect -1 31 0 35
<< ndcontact >>
rect -16 -7 -12 -3
rect 0 -7 4 -3
<< pdcontact >>
rect -16 31 -12 35
rect -8 31 -4 35
rect 0 31 4 35
<< psubstratepcontact >>
rect -18 -15 -14 -11
rect 2 -15 6 -11
<< nsubstratencontact >>
rect -18 39 -14 43
rect 2 39 6 43
<< polysilicon >>
rect -11 35 -9 37
rect -3 35 -1 37
rect -11 -3 -9 31
rect -3 -3 -1 31
rect -11 -9 -9 -7
rect -3 -9 -1 -7
<< polycontact >>
rect -15 22 -11 26
rect -1 13 3 17
<< metal1 >>
rect -21 43 9 44
rect -21 39 -18 43
rect -14 39 2 43
rect 6 39 9 43
rect -21 38 9 39
rect -16 35 -12 38
rect 0 35 4 38
rect -8 7 -4 31
rect -8 3 4 7
rect 0 -3 4 3
rect -16 -10 -12 -7
rect -21 -11 9 -10
rect -21 -15 -18 -11
rect -14 -15 2 -11
rect 6 -15 9 -11
rect -21 -16 9 -15
<< labels >>
rlabel polycontact 1 15 1 15 1 B
rlabel metal1 2 5 2 5 1 Z
rlabel nsubstratencontact -16 41 -16 41 1 +VDD
rlabel nsubstratencontact 4 41 4 41 1 +VDD
rlabel psubstratepcontact -16 -13 -16 -13 1 GND
rlabel psubstratepcontact 4 -13 4 -13 1 GND
rlabel polycontact -13 24 -13 24 1 A
<< end >>
