magic
tech scmos
timestamp 1460491727
<< nwell >>
rect -25 13 13 47
<< pwell >>
rect -25 -36 13 -8
<< ntransistor >>
rect -11 -25 -9 -21
rect -3 -25 -1 -21
<< ptransistor >>
rect -11 31 -9 35
rect -3 31 -1 35
<< ndiffusion >>
rect -12 -25 -11 -21
rect -9 -25 -3 -21
rect -1 -25 0 -21
<< pdiffusion >>
rect -12 31 -11 35
rect -9 31 -8 35
rect -4 31 -3 35
rect -1 31 0 35
<< ndcontact >>
rect -16 -25 -12 -21
rect 0 -25 4 -21
<< pdcontact >>
rect -16 31 -12 35
rect -8 31 -4 35
rect 0 31 4 35
<< psubstratepcontact >>
rect -18 -33 -14 -29
rect 2 -33 6 -29
<< nsubstratencontact >>
rect -18 39 -14 43
rect 2 39 6 43
<< polysilicon >>
rect -11 35 -9 37
rect -3 35 -1 37
rect -11 -21 -9 31
rect -3 -21 -1 31
rect -11 -27 -9 -25
rect -3 -27 -1 -25
<< polycontact >>
rect -15 5 -11 9
rect -1 5 3 9
<< metal1 >>
rect -21 43 9 44
rect -21 39 -18 43
rect -14 39 2 43
rect 6 39 9 43
rect -21 38 9 39
rect -16 35 -12 38
rect 0 35 4 38
rect -8 -11 -4 31
rect -8 -15 4 -11
rect 0 -21 4 -15
rect -16 -28 -12 -25
rect -21 -29 9 -28
rect -21 -33 -18 -29
rect -14 -33 2 -29
rect 6 -33 9 -29
rect -21 -34 9 -33
<< labels >>
rlabel nsubstratencontact -16 41 -16 41 1 +VDD
rlabel nsubstratencontact 4 41 4 41 1 +VDD
rlabel metal1 2 -13 2 -13 1 Z
rlabel psubstratepcontact -16 -31 -16 -31 1 GND
rlabel psubstratepcontact 4 -31 4 -31 1 GND
rlabel polycontact -13 7 -13 7 1 A
rlabel polycontact 1 7 1 7 1 B
<< end >>
