magic
tech scmos
timestamp 1460241092
use NAND2X2  NAND2X2_5
timestamp 1460241041
transform 1 0 -45 0 -1 68
box -25 -18 13 47
use NAND2X2  NAND2X2_3
timestamp 1460241041
transform 1 0 -20 0 -1 68
box -25 -18 13 47
use NAND2X2  NAND2X2_4
timestamp 1460241041
transform 1 0 5 0 -1 68
box -25 -18 13 47
use NAND2X2  NAND2X2_2
timestamp 1460241041
transform 1 0 -45 0 1 -14
box -25 -18 13 47
use NAND2X2  NAND2X2_0
timestamp 1460241041
transform 1 0 -20 0 1 -14
box -25 -18 13 47
use NAND2X2  NAND2X2_1
timestamp 1460241041
transform 1 0 5 0 1 -14
box -25 -18 13 47
use NAND2X2  NAND2X2_6
timestamp 1460241041
transform 1 0 -45 0 -1 -34
box -25 -18 13 47
use NAND2X2  NAND2X2_7
timestamp 1460241041
transform 1 0 -20 0 -1 -34
box -25 -18 13 47
use NAND2X2  NAND2X2_8
timestamp 1460241041
transform 1 0 5 0 -1 -34
box -25 -18 13 47
<< end >>
